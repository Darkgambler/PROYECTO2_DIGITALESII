module synt_glenda( output reg kuka );
   synt_lorita
     synt_perrito
   
